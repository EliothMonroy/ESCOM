library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

entity DIST_RAM is
	GENERIC( 
		NBITS_ADDR : INTEGER := 4;
		NBITS_DATA : INTEGER := 12
		);
    Port ( CLK 	: in  STD_LOGIC;
			  CLR 	: in  STD_LOGIC;
           WE 		: in  STD_LOGIC;
           ADDR 	: in  STD_LOGIC_VECTOR (NBITS_ADDR-1 downto 0);
           DIN 	: in  STD_LOGIC_VECTOR (NBITS_DATA-1 downto 0);
           DOUT 	: out STD_LOGIC_VECTOR (NBITS_DATA-1 downto 0)
			 );
end DIST_RAM;

architecture SINGLE of DIST_RAM is
TYPE MEM_TYPE IS ARRAY ((2**NBITS_ADDR)-1 DOWNTO 0) OF STD_LOGIC_VECTOR(DIN'RANGE);
SIGNAL MEM : MEM_TYPE;
begin
-- ESCRITURA DE MEMORIA
	PMEM : PROCESS( CLK, CLR )
	BEGIN
		IF( CLR = '1' )THEN
			MEM <= (OTHERS => (OTHERS => '0'));
		ELSIF( RISING_EDGE(CLK) )THEN
			IF( WE = '1' )THEN
				MEM(CONV_INTEGER(ADDR)) <= DIN;
			END IF;
		END IF;
	END PROCESS PMEM;
-- LECTURA DE MEMORIA
	DOUT <= MEM(CONV_INTEGER(ADDR));
end SINGLE;