library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity CONT_DECO is
    Port ( CLK : in  STD_LOGIC;
           CLR : in  STD_LOGIC;
           DISPLAY : out  STD_LOGIC_VECTOR (6 downto 0));
end CONT_DECO;

architecture PROGRAMA of CONT_DECO is					-- ABCDEFG
CONSTANT DIGITO0 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0000001";
CONSTANT DIGITO1 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "1001111";
CONSTANT DIGITO2 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0010010";
CONSTANT DIGITO3 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0000110";
CONSTANT DIGITO4 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "1001100";
CONSTANT DIGITO5 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0100100";
CONSTANT DIGITO6 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0100000";
CONSTANT DIGITO7 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0001111";
CONSTANT DIGITO8 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "1111111";
CONSTANT DIGITO9 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0001100";
CONSTANT DIGITOA : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0001000";
CONSTANT DIGITOB : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "1100000";
CONSTANT DIGITOC : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0110001";
CONSTANT DIGITOD : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0000001";
CONSTANT DIGITOE : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0000001";
CONSTANT DIGITOF : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0000001";
SIGNAL Q: STD_LOGIC_VECTOR( 3 DOWNTO 0);
--SIGNAL QDIV: STD_LOGIC_VECTOR( 25 DOWNTO 0);
--SIGNAL QDIV: INTEGER RANGE 0 TO 50000000-1;
--SIGNAL CLK : STD_LOGIC;
begin

----	PDIVISOR : PROCESS( OSC_CLK, CLR )
----	BEGIN
----		IF( CLR = '1' )THEN
----			QDIV <= 0;
----			CLK <= '0';
----		ELSIF( RISING_EDGE( OSC_CLK ) ) THEN
----			QDIV <= QDIV + 1;
----			IF( QDIV = 3 )THEN
----				CLK <= NOT CLK;
----				QDIV <= 0;
----			END IF;
----		END IF;
----	END PROCESS PDIVISOR;
	
	PCONT : PROCESS( CLK, CLR )
	BEGIN
		IF( CLR = '1' )THEN
			Q <= (OTHERS => '0');
		ELSIF( RISING_EDGE( CLK ) ) THEN
			Q <= Q + 1;
		END IF;
	END PROCESS PCONT;
	
	DISPLAY <= 
		DIGITO0 WHEN ( Q <= X"0" ) ELSE
		DIGITO1 WHEN ( Q <= X"1" ) ELSE
		DIGITO2 WHEN ( Q <= X"2" ) ELSE
		DIGITO3 WHEN ( Q <= X"3" ) ELSE
		DIGITO4 WHEN ( Q <= X"4" ) ELSE
		DIGITO5 WHEN ( Q <= X"5" ) ELSE
		DIGITO6 WHEN ( Q <= X"6" ) ELSE
		DIGITO7 WHEN ( Q <= X"7" ) ELSE
		DIGITO8 WHEN ( Q <= X"8" ) ELSE
		DIGITO9 WHEN ( Q <= X"9" ) ELSE
		DIGITOA WHEN ( Q <= X"A" ) ELSE
		DIGITOB WHEN ( Q <= X"B" ) ELSE
		DIGITOC WHEN ( Q <= X"C" ) ELSE
		DIGITOD WHEN ( Q <= X"D" ) ELSE
		DIGITOE WHEN ( Q <= X"E" ) ELSE
		DIGITOF;			
	

end PROGRAMA;

