LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_UNSIGNED.ALL;
USE ieee.std_logic_ARITH.ALL;
USE WORK.PAQUETE.ALL;

entity ROM is
   PORT( ADDRESS : IN  STD_LOGIC_VECTOR( ADDR_N-1 DOWNTO 0);
			  DATA : OUT STD_LOGIC_VECTOR( DATA_N-1 DOWNTO 0)
			  );
end ROM;

ARCHITECTURE PROGRAMA OF ROM IS
signal MROM : MEMORIA := LLENAR_ROM("DATOS.TXT");
BEGIN
	MEMP : PROCESS( ADDRESS )
	BEGIN
		DATA <= MROM( CONV_INTEGER(ADDRESS) );
	END PROCESS MEMP;
END PROGRAMA;