library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

entity DIST_RAM is
	GENERIC( 
		NBITS_ADDR : INTEGER := 4;
		NBITS_DATA : INTEGER := 12
		);
    Port ( CLK 		: in  STD_LOGIC;
           WE 			: in  STD_LOGIC;
           ADDR_WR 	: in  STD_LOGIC_VECTOR (NBITS_ADDR-1 downto 0);
			  ADDR_RD1 	: in  STD_LOGIC_VECTOR (NBITS_ADDR-1 downto 0);
			  ADDR_RD2 	: in  STD_LOGIC_VECTOR (NBITS_ADDR-1 downto 0);
           DIN 		: in  STD_LOGIC_VECTOR (NBITS_DATA-1 downto 0);
           DOUT1 		: out STD_LOGIC_VECTOR (NBITS_DATA-1 downto 0);
			  DOUT2 		: out STD_LOGIC_VECTOR (NBITS_DATA-1 downto 0)
			  );
end DIST_RAM;

architecture DUAL of DIST_RAM is
TYPE MEM_TYPE IS ARRAY ((2**NBITS_ADDR)-1 DOWNTO 0) OF STD_LOGIC_VECTOR(DIN'RANGE);
SIGNAL MEM : MEM_TYPE;

begin
-- ESCRITURA DE MEMORIA
	PMEM : PROCESS( CLK )
	BEGIN
		IF( RISING_EDGE(CLK) )THEN
			IF( WE = '1' )THEN
				MEM(CONV_INTEGER(ADDR_WR)) <= DIN;
			END IF;
		END IF;
	END PROCESS PMEM;
-- LECTURA DE MEMORIA
	DOUT1 <= MEM(CONV_INTEGER(ADDR_RD1));
	DOUT2 <= MEM(CONV_INTEGER(ADDR_RD2));
end DUAL;

