library ieee;
use ieee.std_logic_1164.all;
library lattice;
use lattice.components.all;
entity ha is
	port(
		A0: in std_logic;
		B0: in std_logic;
		S0: out std_logic;
		c0: out std_logic);
end ha;
architecture ha0 of ha is
begin
	
end;