LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY CONT_GEN IS
	PORT(																					
		CLK, CLR : IN STD_LOGIC;
		D : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		OPER : IN STD_LOGIC_VECTOR( 1 DOWNTO 0 );
		Q : INOUT STD_LOGIC_VECTOR( 7 DOWNTO 0 )
	); 
END CONT_GEN;

ARCHITECTURE ACONT OF CONT_GEN IS
BEGIN
	PCONT : PROCESS( CLK, CLR )
	BEGIN		
		IF( CLR = '1' )THEN
			Q <= (OTHERS => '0');
		ELSIF( CLK'EVENT AND CLK = '1' )THEN
			CASE OPER IS
				WHEN "00" => 
					Q <= D;
				WHEN "01" => 
					Q <= Q;	
				WHEN "10" =>
					Q <= Q + 1;
				WHEN OTHERS => 
					Q <= Q - 1;
			END CASE;
		END IF;
	END PROCESS PCONT;
END ACONT;

