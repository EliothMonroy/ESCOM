library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity Decodificador is

port( 
	a: in std_logic_vector ( 5 downto 0 );
	s: out std_logic_vector ( 15 downto 0 ) );
	attribute loc: string;
	attribute loc of a:signal is "p4,p5,p6,p7,p8,9";
	attribute loc of s:signal is "p111,p112,p113,p114,p115,p116,p120,p121,p122,p123,p124,p125,p130,p131,p132,p133";

end;

architecture dec of Decodificador is
begin
	process(a) begin
		case a is--Catodo (Prende con unos)
		         --             "123456789ABCDEFG"
			when "000000" =>s<= "1111111101100000";--0
			when "000001" =>s<= "0011000000000000";--1
			when "000010" =>s<= "1110111000001100";--2
			when "000011" =>s<= "1111110000001100";--3
			when "000100" =>s<= "0011000100001100";--4
			when "000101" =>s<= "1101110100001100";--5
			when "000110" =>s<= "1101111100001100";--6
			when "000111" =>s<= "1111000000000000";--7
			when "001000" =>s<= "1111111100001100";--8
			when "001001" =>s<= "1111000100001100";--9
		         --             "123456789ABCDEFG"
			when "001010" =>s<= "1111001100001100";--A(10)
			when "001011" =>s<= "0001111100001100";--b(11)
			when "001100" =>s<= "1100111100000000";--C(12)
			when "001101" =>s<= "0011111000001100";--d(13)
			when "001110" =>s<= "1100111100001100";--E(14)
			when "001111" =>s<= "1100001100001100";--F(15)
			when "010000" =>s<= "1101111100000100";--G(16)
			when "010001" =>s<= "0011001100001100";--H(17)
			when "010010" =>s<= "1100110000000011";--I(18)
			when "010011" =>s<= "1100010000000011";--J(19)
			when "010100" =>s<= "0000000001010011";--k(20)
		         --             "123456789ABCDEFG"
			when "010101" =>s<= "0000111100000000";--L(21)
			when "010110" =>s<= "0011001111000000";--M(22)
			when "010111" =>s<= "0011001110010000";--N(23)
			when "011000" =>s<= "1111111100000000";--O(24)
			when "011001" =>s<= "1110001100001100";--P(25)
			when "011010" =>s<= "1111111100010000";--Q(26)
			when "011011" =>s<= "1110001100011100";--R(27)
			when "011100" =>s<= "1000010100001001";--s(28)
			when "011101" =>s<= "1100000000000011";--T(29)
			when "011110" =>s<= "0011111100000000";--U(30)
		         --             "123456789ABCDEFG"
			when "011111" =>s<= "0000000011000000";--V(31)
			when "100000" =>s<= "0011001100110000";--W(32)
			when "100001" =>s<= "0000000011110000";--X(33)
			when "100010" =>s<= "0000000011000001";--Y(34)
			when "100011" =>s<= "1100110001100000";--Z(35)
			when others   =>s<= "1111111111111111";
		end case;
	end process ; -- process
end dec;

